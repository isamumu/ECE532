// DCT module to compute the Discrete Cosine Transform
module DCT(
#(
  parameter PICTURE_SIZE = 32
)
(

);

endmodule

module compute_am(input l, );

endmodule 